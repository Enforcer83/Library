*---------- DMN2990UFA Spice Model ----------

*NMOS
.SUBCKT DMN2990UFA 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1E-006  W = 1E-006 
RD 10 1 0.3743 
RS 30 3 0.001 
RG 20 2 113 
CGS 2 3 2.5E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1  VFB 1 
CGD 13 14 8E-011 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 3 10  DSUB 
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1E+006  ETA = 0.01  VTO = 0.8716 
+ TOX = 6E-008  NSUB = 1.886E+016  KP = 2.108  U0 = 400  KAPPA = 10.7 
.MODEL DCGD D  CJO = 1.594E-011  VJ = 0.2646  M = 0.429 
.MODEL DSUB D  IS = 2.265E-009  N = 1.422  RS = 1.834  BV = 25  CJO = 2.7E-012  VJ = 0.2048  M = 0.1841 
.MODEL DLIM D  IS = 0.0001 
.ENDS


*Diodes DMN2990UFA Spice Model v1.0 Last Revised 2012/11/30