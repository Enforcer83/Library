* ADG658 MACROMODEL MODEL CAN ONLY RUN ON SPICE2
* Description: Converter
* Generic Desc: 3V/5V  4/8 Channel Analog muxs
* Developed by: Y.WONG
* Revision History: 08/10/2012 - Updated to new header style
* 1.1 (11/2008)
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
*
* END Notes
*
* Connections
*      1  = S5
*      2  = S7
*      3  = D
*      4  = S8
*      5  = S6
*      6  = /EN
*      7  = VSS
*      8  = GND
*      9  = A2
*      10 = A1
*      11 = A0
*      12 = S4
*      13 = S1
*      14 = S2
*      15 = S3
*      16 = VDD
*****************
.SUBCKT ADG658 S5 S7 D S8 S6 NEN VSS GND A2 A1 A0 S4 S1 S2 S3 VDD
RL1 VDD GND 5000MEG
RL2 VSS GND 5000MEG
CEN NEN GND 2p
CA0 A2 GND 2p
CA1 A1 GND 2p
CA2 A2 GND 2p
DENA NEN VDD DY
DENB VSS NEN DY
DA0A A0 VDD DY
DA0B VSS A0 DY
DA1A A1 VDD DY
DA1B VSS A1 DY
DA2A A2 VDD DY
DA2B VSS A2 DY
X9 NEN A0 A1 A2 VDD GND 17 18 19 20 21 22 23 24 DECODER
X1 S1 D 17 VDD GND VSS NEN  HIGHONSWITCH
X2 S2 D 18 VDD GND VSS NEN  HIGHONSWITCH
X3 S3 D 19 VDD GND VSS NEN  HIGHONSWITCH
X4 S4 D 20 VDD GND VSS NEN  HIGHONSWITCH
X5 S5 D 21 VDD GND VSS NEN  HIGHONSWITCH
X6 S6 D 22 VDD GND VSS NEN  HIGHONSWITCH
X7 S7 D 23 VDD GND VSS NEN  HIGHONSWITCH
X8 S8 D 24 VDD GND VSS NEN  HIGHONSWITCH
CS12 S1 S2 0.01p
CS13 S1 S3 0.01p
CS14 S1 S4 0.01p
CS15 S1 S5 0.01p
CS16 S1 S6 0.01p
CS17 S1 S7 0.01p
CS18 S1 S8 0.01p
CS23 S2 S3 0.01p
CS24 S2 S4 0.01p
CS25 S2 S5 0.01p
CS26 S2 S6 0.01p
CS27 S2 S7 0.01p
CS28 S2 S8 0.01p
CS34 S3 S4 0.01p
CS35 S3 S5 0.01p
CS36 S3 S6 0.01p
CS37 S3 S7 0.01p
CS38 S3 S8 0.01p
CS45 S4 S5 0.01p
CS46 S4 S6 0.01p
CS47 S4 S7 0.01p
CS48 S4 S8 0.01p
CS56 S5 S6 0.01p
CS57 S5 S7 0.01p
CS58 S5 S8 0.01p
CS67 S6 S7 0.01p
CS68 S6 S8 0.01p
CS78 S7 S8 0.01p
*MODELS USED
.MODEL DY D(IS=1E-14 N=0.04 RS=30)
.ENDS

*****************
* 3 to 8 with Enable Low Decoder
*
* Connections
*      101 = /EN
*      102 = A0
*      103 = A1
*      104 = A2
*      105 = VDD
*      106 = GND
*      107 = D1
*      108 = D2
*      109 = D3
*      110 = D4
*      111 = D5
*      112 = D6
*      113 = D7
*      114 = D8
*****************

.SUBCKT DECODER 101 102 103 104 105 106 107 108 109 110 111 112 113 114
SEN 150 106 101 106 SMOD2
SA0 115 106 102 106 SMOD2
SA1 116 106 103 106 SMOD2
SA2 117 106 104 106 SMOD2
SD1A 105 118 150 106 SMOD2
SD1B 118 119 115 106 SMOD2
SD1C 119 120 116 106 SMOD2
SD1D 120 121 117 106 SMOD2
SD2A 105 122 150 106 SMOD2
SD2B 122 123 102 106 SMOD2
SD2C 123 124 116 106 SMOD2
SD2D 124 125 117 106 SMOD2
SD3A 105 126 150 106 SMOD2
SD3B 126 127 115 106 SMOD2
SD3C 127 128 103 106 SMOD2
SD3D 128 129 117 106 SMOD2
SD4A 105 130 150 106 SMOD2
SD4B 130 131 102 106 SMOD2
SD4C 131 132 103 106 SMOD2
SD4D 132 133 117 106 SMOD2
SD5A 105 134 150 106 SMOD2
SD5B 134 135 115 106 SMOD2
SD5C 135 136 116 106 SMOD2
SD5D 136 137 104 106 SMOD2
SD6A 105 138 150 106 SMOD2
SD6B 138 139 102 106 SMOD2
SD6C 139 140 116 106 SMOD2
SD6D 140 141 104 106 SMOD2
SD7A 105 142 150 106 SMOD2
SD7B 142 143 115 106 SMOD2
SD7C 143 144 103 106 SMOD2
SD7D 144 145 104 106 SMOD2
SD8A 105 146 150 106 SMOD2
SD8B 146 147 102 106 SMOD2
SD8C 147 148 103 106 SMOD2
SD8D 148 149 104 106 SMOD2
REN 150 105 5G
RA0 115 105 5G
RA1 116 105 5G
RA2 117 105 5G
RD1 121 106 5G
RD2 125 106 5G
RD3 129 106 5G
RD4 133 106 5G
RD5 137 106 5G
RD6 141 106 5G
RD7 145 106 5G
RD8 149 106 5G
ED1 107 106 121 106 1
ED2 108 106 125 106 1
ED3 109 106 129 106 1
ED4 110 106 133 106 1
ED5 111 106 137 106 1
ED6 112 106 141 106 1
ED7 113 106 145 106 1
ED8 114 106 149 106 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-03 ROFF=1E11 VON=2.0 VOFF=0.8)
.ENDS

****************
* Logic High On Switch
*
* Connections
*      101 = S
*      102 = D
*      103 = VIN
*      104 = VDD
*      105 = GND
*      106 = VSS
*      107 = /EN
*****************

.SUBCKT HIGHONSWITCH  101 102 103 104 105 106 107

x1 103 104 105 108 BUFF
X2 108 109 104 106 105 VSENSE
X3 109 110 107 105 ENABLE
X4 110 105 111 ENABLEDELAY
X5 101 102 111 104 105 106 SWITCH

*MODELS USED
.ENDS

****************
* Switch
*
* Connections
*      201 = S
*      202 = D
*      203 = VIN
*      204 = VDD
*      205 = GND
*      206 = VSS
*****************

.SUBCKT SWITCH  201 202 203 204 205 206

*ANALOG SWITCH
EBuffer 214 205 202 205 1
S1 210 202 203 205 SMOD1
Vo2 214 219 0
EVDD 219 220 204 205 1
SN 210 209 205 220 SMOD7
Vo1 205 218 0
EVSS 217 218 206 205 1
SP 210 208 214 217 SMOD8
Xn 215 209 214 205 204 206 VCRN
Xp 207 208 214 205 204 206 VCRP
RS1 201 207 1
RS2 201 215 1

DS1 201 204 DX
DS2 206 201 DX
DD1 202 204 DX
DD2 206 202 DX

*ON OFF ISOLATION*
CSD 201 202 0.201p

*BANDWIDTH *
CSB 201 206 2.1p
CDB 202 204 2.1p

*CHARGE INJECTION
CGS 201 203 0.167p
CGD 202 203 0.167p

*MODELS USED
.MODEL SMOD1 VSWITCH(RON=1 ROFF=7E11 VON=2.0 VOFF=0.8)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.81 VOFF=0.79)
.MODEL SMOD8 VSWITCH(RON=1E-3 ROFF=1E11 VON=1.21 VOFF=1.19)
.MODEL DX D(IS=1E-12 N=0.04 RS=120)
.ENDS

*****************
* BUFF LOGIC
*
* Connections
*      201 = INPUT
*      202 = VDD
*      203 = GND
*      204 = OUTPUT
*****************
.SUBCKT BUFF 201 202 203 204
SBUFF 205 203 201 203 SMOD2
RBUFF 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* ENABLE DELAY
*
* Connections
*      301 = INPUT
*      302 = COM
*      303 = OUTPUT
*****************
.SUBCKT ENABLEDELAY 301 302 303

EENBUFFER 304 302 301 302 1
RFEN 304 306 45k
CFEN 306 302 5p
DBREAKEN 306 305 DZ
RBEN 305 304 17k
EENBUFFEROUT 303 302 306 302 1

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* Enable ON/OFF
*
* Connections
*      501 = INPUT
*      502 = OUTPUT
*      503 = VIN
*      504 = GND
*****************
.SUBCKT ENABLE 501 502 503 504
SENABLE 501 505 503 504 SMOD2
RD0 505 504 5G
EBUFFER 502 504 505 504 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* OPERATING VOLTAGE
*
* Connections
*      601 = INPUT
*      602 = OUTPUT
*      603 = VDD
*      604 = VSS
*      605 = GND
*****************
.SUBCKT VSENSE 601 602 603 604 605
SD1 601 606 603 605 SMOD3
SD2 606 607 603 605 SMOD4
SD3 607 608 605 604 SMOD5
SD4 608 609 605 604 SMOD6
SD5 609 602 603 604 SMOD7
RD0 602 605 5G

*MODELS USED
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E11 VON=2 VOFF=1.9)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)
.MODEL SMOD5 VSWITCH(RON=1E-3 ROFF=1E11 VON=0 VOFF=-0.1)
.MODEL SMOD6 VSWITCH(RON=1E-3 ROFF=1E11 VON=6 VOFF=6.1)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)

.ENDS

*****************
* Voltage Controlled Resistance n-channel
*
* Connections
*      701 = R+
*      702 = R-
*      704 = V+
*      705 = V-
*      707 = VDD
*      711 = VSS
*****************
.SUBCKT VCRN 701 702 704 705 707 711
vtn 708 0 0.8
ERES 701 703 VALUE={285*V(706,0)*(1/(V(707,0)-V(704,705)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS

*****************
* Voltage Controlled Resistance p-channel
*
* Connections
*      701 = R+
*      702 = R-
*      704 = V+
*      705 = V-
*      707 = VDD
*      711 = VSS
*****************
.SUBCKT VCRP 701 702 704 705 707 711
vtp 708 0 1.2
ERES 701 703 VALUE={246*V(706,0)*(1/(V(704,705)-V(711,0)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS




