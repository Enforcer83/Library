*BEGIN MODEL LMH6609
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
* For more information, and our latest models,
* please visit the models section of our website at
*       http://www.national.com/models/
*////////////////////////////////////////////////////////////////////
*MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THRU
*THE SUPPLY RAILS, GAIN AND PHASE, SLEW RATE, COMMON MODE
*REJECTION, POWER SUPPLY REJECTION ON BOTH RAILS, INPUT
*VOLTAGE NOISE WITH 1/F,INPUT CURRENT NOISE WITH 1/F,
*OUPUT IMPEDANCE, INPUT CAPACITANCE, INPUT BIAS CURRENT,
*INPUT COMMON MODE RANGE,INPUT OFFSET, HIGH CLOAD DRIVE
*CAPABILITY, OUTPUT CLAMPS TO THE RAIL, AND QUIESCENT
*SUPPLY CURRENT.

*MODEL TEMP RANGE IS -40 TO +85 DEG C.
*///////////////////////////////////////////////////////
**********************************
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   4   5  2  1
.SUBCKT LMH6609 3 4 5 2 1
* BEGIN MODEL PROGRAMMING
* USE +- 5 VOLT GROUP OR +-3.3 V GROUP BY
* UNCOMMENTING DESIRED GROUP (3 LINES)
* FOR SUPPLY VALUES BETWEEN +-3.3 AND +-5
* LINEARLY INTERPOLATE VALUES
************
* BEGIN +-5 VOLT GROUP
************
* R68 AND R69 MODIFY VOLTAGE NOISE
* G5 MODIFIES BANDWIDTH AND SLEW
R68 27 51 17
R69 52 50 17
G5 39 0 42 43 -1E-3
* END +-5 VOLT GROUP
************
* BEGIN +-3.3 VOLT GROUP
************
* R68 AND R69 MODIFY VOLTAGE NOISE
* G5 MODIFIES BANDWIDTH AND SLEW
*R68 27 51 125
*R69 52 50 125
*G5 39 0 42 43 -0.85E-3
* END +-3.3 VOLT GROUP
* END MODEL PROGRAMMING
Q17 2 6 7 QOP
Q21 5 8 7 QON
D5 1 5 DD
D6 2 1 DD
D7 9 0 DIN
D8 10 0 DIN
I8 0 9 0.1E-3
I9 0 10 0.1E-3
E2 11 0 2 0 1
E3 12 0 5 0 1
D9 13 0 DVN
D10 14 0 DVN
I10 0 13 2E-3
I11 0 14 2E-3
E4 15 4 13 14 1
G2 3 15 9 10 0.45E-4
R22 2 5 66E3
E5 16 0 12 0 1
E6 17 0 11 0 1
E7 18 0 19 0 1
R30 16 20 1E3
R31 17 21 1E3
R32 18 22 1E3
R33 0 20 0.1
R34 0 21 0.1
R35 0 22 0.1
E10 23 3 22 0 0.63
R36 24 19 1E3
R37 19 25 1E3
C6 16 20 1000E-12
C7 17 21 2000E-12
C8 18 22 2000E-12
E11 26 23 21 0 0.63
E12 27 26 20 0 0.91
Q22 11 28 8 QDP
Q23 12 28 6 QDN
I12 5 2 -3.7E-3
I13 12 8 0.6E-3
I14 6 11 0.6E-3
R38 0 29 10
R39 0 28 10
C9 29 0 15E-12
C10 28 0 12E-12
E15 30 31 32 0 1
E16 31 33 32 0 1
E17 34 0 31 0 1
D11 35 12 DD
D12 11 36 DD
V11 33 36 1.75
V12 35 30 1.75
I15 0 37 1E-3
D13 37 0 DD
V13 32 37 -0.6551
C11 31 0 2.9E-12
D14 38 39 DD
D15 39 40 DD
R40 39 31 5
R41 0 39 600E3
C12 15 0 1.2E-12
C13 27 0 1.2E-12
R43 7 41 7
G3 29 0 31 0 0.1
G4 28 0 29 0 0.1
L1 41 1 4E-9
R45 41 1 100
E20 38 34 32 0 1
E21 40 34 32 0 -1
C15 15 27 0.2E-12
R49 44 45 210
R50 44 46 210
I16 12 47 3.1E-3
R51 42 48 1527
R52 43 48 1527
V14 44 49 0.7
V15 12 48 0
C17 42 43 0.02E-12
D18 50 12 DIC
D19 51 12 DIC
E25 25 0 3 0 1
E26 24 0 15 0 1
C18 1 0 0.1E-12
R58 31 30 1E9
R59 33 31 1E9
R60 4 15 1E9
R61 3 23 1E9
R62 23 26 1E9
R63 26 27 1E9
V16 15 50 0.57E-3
R64 34 40 1E9
R65 34 38 1E9
Q28 42 52 45 QIN
Q29 43 51 46 QIN
Q30 49 47 11 QIN
Q31 47 47 11 QIN
G6 5 2 5 2 1E-3
I17 0 50 5.2E-6
I18 0 51 5.2E-6
R70 0 32 1E9
.MODEL QDP PNP
.MODEL QDN NPN
.MODEL QON NPN VAF=150 BF=200 IKF=1.5 RE=1 RC=9
.MODEL QOP PNP VAF=150 BF=200 IKF=1.5 RE=1 RC=9
.MODEL QIN NPN VAF=150 BF=320 IKF=0.005 RE=1 RC=1
.MODEL DD D
.MODEL DVN D KF=1E-14
.MODEL DIN D KF=26E-14
.MODEL DIC D RS=500
.ENDS
*END MODEL LMH6609